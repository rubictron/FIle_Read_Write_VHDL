-- No default header stored in vhdlConfig.txt
entity top_level is
   port (

   );
end entity rtl_BLOCKNAME;

architecture rtl of rtl_BLOCKNAME is

begin

end architecture rtl;library ieee;
use ieee.std_logic_1164.all;